module bram(
    input wire clk,
    input wire rst,
    output wire data
);
endmodule