`define INST_BURST_NUM 8'h7