`define INST_BURST_NUM 8'h7
`define DATA_BURST_NUM 8'h7